package adder_testbench_pkg;
  import uvm_pkg::*;
  
  // Include files here
  
endpackage
