interface switch_input_interface(input clk);
  
	//Define the input interface signals

	//Define the driver clocking block

	//Define the driver modport

	//Define the monitor clocking block 

	//Define the monitor modport  


endinterface

