package switch_testbench_pkg;
  import uvm_pkg::*;
  
  `include "switch_sequence.sv"
  `include "switch_driver.sv"
  `include "switch_monitor_input.sv"
  `include "switch_monitor_output.sv"
  `include "switch_scoreboard.sv"
  `include "switch_agent_input.sv"
  `include "switch_agent_output.sv"
  `include "switch_env.sv"
  `include "switch_test.sv"

endpackage
  
