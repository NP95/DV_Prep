interface adder_interface();
  
  //Define the interface ports below

endinterface
