package phases_testbench_pkg;
  import uvm_pkg::*;
  
  `include "uvm_cmpt_2.sv"
  `include "uvm_cmpt_1.sv"
  `include "uvm_test_1.sv"

endpackage
  
