interface switch_output_interface(input clk);
  
	//Define output interface signals

	//Define the clocking block

	//Define the modport

endinterface
