interface ram_interface(input clk);
  
  logic [7:0] address;
  wire logic [15:0] data;
  logic rd_req;
  logic wr_req;
  logic rd_valid;

  //Add driver clocking block

  //Define driver modport

  //Add monitor clocking block

  //Define monitor modport
  
endinterface
