package reporting_testbench_pkg;
  import uvm_pkg::*;
  
  `include "uvm_reporting.sv"
  `include "uvm_test_1.sv"

endpackage
  
