  `include "adder_sequence_item.sv"
  `include "adder_driver.sv"
  `include "adder_monitor.sv"
  `include "adder_env.sv"
